`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// 
// Module Name: SignExtend
// 
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module SignExtend(in, out);

    input [4:0] in;
    
    output reg [31:0] out;
    
    always @(in) begin
        out = in;
    end
