`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Lab D2L group 38, bench 28 
//Team Members: Christopher Hughes, Sarah Wiltbank
//Percent Effort: Christopher 50/50 Sarah
//
// ECE369A - Computer Architecture
// Laboratory  
// Module - PCAdder.v
// Description - 32-Bit program counter (PC) adder.
// 
// INPUTS:-
// PCResult: 32-Bit input port.
// 
// OUTPUTS:-
// PCAddResult: 32-Bit output port.
//
// FUNCTIONALITY:-
// Design an incrementor (or a hard-wired ADD ALU whose first input is from the 
// PC, and whose second input is a hard-wired 4) that computes the current 
// PC + 4. The result should always be an increment of the signal 'PCResult' by 
// 4 (i.e., PCAddResult = PCResult + 4).
////////////////////////////////////////////////////////////////////////////////

module PCAdder(PCResult, PCAddResult);

    input [31:0] PCResult;


    output  reg [31:0] PCAddResult;

   initial begin
        PCAddResult <= 0;
    end
    
    
      always @(*) begin
        
           PCAddResult <= PCResult + 4;
        
      end

endmodule
